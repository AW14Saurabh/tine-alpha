LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY tine_alpha;

PACKAGE fetch_stage_const IS

    CONSTANT NOP_INST : STD_LOGIC_VECTOR(7 DOWNTO 0) := x"00";

END fetch_stage_const;