LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE alu_const IS

    CONSTANT AO_SKNV : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    CONSTANT AO_SKIP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
    CONSTANT AO_SKNE : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
    CONSTANT AO_SKE : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
    CONSTANT AO_SKL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
    CONSTANT AO_SKLE : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
    CONSTANT AO_SKG : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
    CONSTANT AO_SKGE : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
    CONSTANT AO_AND : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
    CONSTANT AO_NOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
    CONSTANT AO_SLL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
    CONSTANT AO_SRL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
    CONSTANT AO_SLU : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";
    CONSTANT AO_SL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";
    CONSTANT AO_SUB : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110";
    CONSTANT AO_ADD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111";

END alu_const;