LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY tine_alpha;

PACKAGE address_stage_const IS

    CONSTANT RST_IP_REG : STD_LOGIC_VECTOR(7 DOWNTO 0) := x"00";

END address_stage_const;